`timescale 1ns / 1ps

module fifo #(parameter DEPTH=8, DWIDTH=16)
    (
            input               	rstn,               // Active low reset
                                    clk,                // Clock
                                    wr_en, 				// Write enable
                                    rd_en, 				// Read enable
            input      [DWIDTH-1:0] din, 				// Data written into FIFO
            output reg [DWIDTH-1:0] dout, 				// Data read from FIFO
            output              	empty, 				// FIFO is empty when high
                                    full 				// FIFO is full when high
    );
    
    
      reg [$clog2(DEPTH)-1:0]   wptr;
      reg [$clog2(DEPTH)-1:0]   rptr;
    
      reg [DWIDTH-1 : 0]    fifo[DEPTH];
    
      always_ff @ (posedge clk) begin
        if (!rstn) begin
          wptr <= 0;
        end else begin
          if (wr_en & !full) begin
            fifo[wptr] <= din;
            wptr <= wptr + 1;
          end
        end
      end
    
    
      always_ff @ (posedge clk) begin
        if (!rstn) begin
          rptr <= 0;
        end else begin
          if (rd_en & !empty) begin
            dout <= fifo[rptr];
            rptr <= rptr + 1;
          end
          else dout = {DWIDTH{1'bx}};
        end
      end
    
      assign full  = (wptr + 1) == rptr;
      assign empty = wptr == rptr;
    endmodule